module gate_not(input a, output out);
    assign out = !a;    
endmodule


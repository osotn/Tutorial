module gate_or(input a, input b, output out);
    assign out = a | b;    
endmodule

